module CPU 